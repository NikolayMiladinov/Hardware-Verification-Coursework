package my_pkg;
`include "transaction.sv"
`include "generator.sv"
`include "gpio_intf.sv"
`include "driver.sv"
`include "environment.sv"
`include "test.sv"
// `include "monitor.sv"
// `include "scoreboard.sv"
endpackage